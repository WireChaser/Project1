// megafunction wizard: %ROM: 2-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram

// ============================================================
// File Name: ram_result.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.0.0 Build 614 04/24/2018 SJ Lite Edition
// ************************************************************


//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions
//and other software and tools, and its AMPP partner logic
//functions, and any output files from any of the foregoing
//(including device programming or simulation files), and any
//associated documentation or information are expressly subject
//to the terms and conditions of the Intel Program License
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.

`timescale 1 ps / 1 ps

module ram_result 
   #(parameter ADDR_WIDTH = 7,
	       RESULT_WIDTH = 24)
   (address_a,
   address_b,
   clock,
   data_a,
   data_b,
   q_a,
   q_b,
   wren_a,
   wren_b);

   input [ADDR_WIDTH-1:0]  address_a, address_b;
   input [RESULT_WIDTH-1:0]  data_a, data_b;
   input clock;
   input logic wren_a, wren_b;
   output[RESULT_WIDTH-1:0]  q_a, q_b;

   altsyncram altsyncram_component (
     		 .address_a (address_a),
                 .address_b (address_b),
     		 .clock0 (clock),
     		 .data_a (data_a),
     		 .data_b (data_b),
     		 .wren_a (wren_a),
     		 .wren_b (wren_b),
     		 .q_a (q_a),
     		 .q_b (q_b)
     		 ,
     		 .aclr0 (),
     		 .aclr1 (),
     		 .addressstall_a (),
     		 .addressstall_b (),
     		 .byteena_a (),
     		 .byteena_b (),
     		 .clock1 (),
     		 .clocken0 (),
     		 .clocken1 (),
     		 .clocken2 (),
     		 .clocken3 (),
     		 .eccstatus (),
      		 .rden_a (),
     		 .rden_b ()
  	   );
   defparam
      altsyncram_component.address_reg_b = "CLOCK0",
      altsyncram_component.clock_enable_input_a = "BYPASS",
      altsyncram_component.clock_enable_input_b = "BYPASS",
      altsyncram_component.clock_enable_output_a = "BYPASS",
      altsyncram_component.clock_enable_output_b = "BYPASS",
      altsyncram_component.indata_reg_b = "CLOCK0",
      altsyncram_component.intended_device_family = "Cyclone V",
      altsyncram_component.lpm_type = "altsyncram",
      altsyncram_component.numwords_a = 2**ADDR_WIDTH,
      altsyncram_component.numwords_b = 2**ADDR_WIDTH,
      altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
      altsyncram_component.outdata_aclr_a = "NONE",
      altsyncram_component.outdata_aclr_b = "NONE",
      altsyncram_component.outdata_reg_a = "UNREGISTERED",
      altsyncram_component.outdata_reg_b = "UNREGISTERED",
      altsyncram_component.power_up_uninitialized = "FALSE",
      altsyncram_component.ram_block_type = "M10K",
      altsyncram_component.widthad_a = ADDR_WIDTH,
      altsyncram_component.widthad_b = ADDR_WIDTH,
      altsyncram_component.width_a = RESULT_WIDTH,
      altsyncram_component.width_b = RESULT_WIDTH,
      altsyncram_component.width_byteena_a = 1,
      altsyncram_component.width_byteena_b = 1,
      altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0";
	
endmodule 
